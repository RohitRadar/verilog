`timescale 1ns/1ps

module djikstras_tb();
	reg clk_50;
	wire [63:0] direction_out;
	reg [7:0] starting_node;
	reg [7:0] ending_node;
	
	integer clk_i,cycle=20;
	djikstras DUT(.clk_50(clk_50),
					  .direction_out(direction_out),
					  .starting_node(starting_node),
					  .ending_node(ending_node)
	);
	initial
	begin
		starting_node=1;
		ending_node=22;
		for(clk_i=0;clk_i<20000;clk_i=clk_i+1)
		begin
			clk_50=1'b0;
			#(cycle/2);
			clk_50=1'b1;
			#(cycle/2);
		end
		starting_node=22;
		ending_node=17;
		for(clk_i=0;clk_i<20000;clk_i=clk_i+1)
		begin
			clk_50=1'b0;
			#(cycle/2);
			clk_50=1'b1;
			#(cycle/2);
		end
		starting_node=17;
		ending_node=3;
		for(clk_i=0;clk_i<20000;clk_i=clk_i+1)
		begin
			clk_50=1'b0;
			#(cycle/2);
			clk_50=1'b1;
			#(cycle/2);
		end
		starting_node=3;
		ending_node=14;
		for(clk_i=0;clk_i<20000;clk_i=clk_i+1)
		begin
			clk_50=1'b0;
			#(cycle/2);
			clk_50=1'b1;
			#(cycle/2);
		end
		starting_node=14;
		ending_node=23;
		for(clk_i=0;clk_i<20000;clk_i=clk_i+1)
		begin
			clk_50=1'b0;
			#(cycle/2);
			clk_50=1'b1;
			#(cycle/2);
		end
		starting_node=23;
		ending_node=30;
		for(clk_i=0;clk_i<20000;clk_i=clk_i+1)
		begin
			clk_50=1'b0;
			#(cycle/2);
			clk_50=1'b1;
			#(cycle/2);
		end
		starting_node=30;
		ending_node=36;
		for(clk_i=0;clk_i<20000;clk_i=clk_i+1)
		begin
			clk_50=1'b0;
			#(cycle/2);
			clk_50=1'b1;
			#(cycle/2);
		end
		starting_node=36;
		ending_node=26;
		for(clk_i=0;clk_i<20000;clk_i=clk_i+1)
		begin
			clk_50=1'b0;
			#(cycle/2);
			clk_50=1'b1;
			#(cycle/2);
		end
		starting_node=26;
		ending_node=32;
		for(clk_i=0;clk_i<20000;clk_i=clk_i+1)
		begin
			clk_50=1'b0;
			#(cycle/2);
			clk_50=1'b1;
			#(cycle/2);
		end
		starting_node=32;
		ending_node=37;
		for(clk_i=0;clk_i<20000;clk_i=clk_i+1)
		begin
			clk_50=1'b0;
			#(cycle/2);
			clk_50=1'b1;
			#(cycle/2);
		end
		starting_node=37;
		ending_node=1;
		for(clk_i=0;clk_i<20000;clk_i=clk_i+1)
		begin
			clk_50=1'b0;
			#(cycle/2);
			clk_50=1'b1;
			#(cycle/2);
		end
		$finish;
	end
endmodule
